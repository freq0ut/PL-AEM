library ieee;
use ieee.std_logic_1164.all;

ENTITY Multiplier_Encoder_7_Bit IS
	PORT(
		A 	: 	IN  std_logic_vector  (6 DOWNTO 0);
		B 	: 	OUT std_logic_vector (10 DOWNTO 0)
	);
END Multiplier_Encoder_7_Bit;

ARCHITECTURE behavioral OF Multiplier_Encoder_7_Bit IS
BEGIN

WITH A SELECT
		B <= 
			-- 11 bit out and 7 bit in
			"00000000000" WHEN "0000000", -- 0
			"00001000000" WHEN "0000001", -- 1
			"00000001000" WHEN "0000010", -- 2
			"00000001001" WHEN "0000011", -- 3

			"00001001001" WHEN "0000100", -- 4
			"00000001010" WHEN "0000101", -- 5
			"00001001010" WHEN "0000110", -- 6
			"00011000000" WHEN "0000111", -- 7

			"00010001010" WHEN "0001000", -- 8
			"00000001011" WHEN "0001001", -- 9
			"00001001011" WHEN "0001010", -- 10
			"00011011000" WHEN "0001011", -- 11

			"00010001011" WHEN "0001100", -- 12
			"00000011010" WHEN "0001101", -- 13
			"00100000001" WHEN "0001110", -- 14
			"00100000000" WHEN "0001111", -- 15

			"00011001011" WHEN "0010000", -- 16
			"00000001100" WHEN "0010001", -- 17
			"00001001100" WHEN "0010010", -- 18
			"00100011000" WHEN "0010011", -- 19

			"00010001100" WHEN "0010100", -- 20
			"00000101010" WHEN "0010101", -- 21
			"00100011001" WHEN "0010110", -- 22
			"00100111000" WHEN "0010111", -- 23

			"00011001100" WHEN "0011000", -- 24
			"00000011011" WHEN "0011001", -- 25
			"00001011011" WHEN "0011010", -- 26
			"00101100000" WHEN "0011011", -- 27

			"00101000010" WHEN "0011100", -- 28
			"00101010000" WHEN "0011101", -- 29
			"00101000001" WHEN "0011110", -- 30
			"00101000000" WHEN "0011111", -- 31

			"00100001100" WHEN "0100000", -- 32
			"00000001101" WHEN "0100001", -- 33
			"00001001101" WHEN "0100010", -- 34
			"00101011000" WHEN "0100011", -- 35

			"00010001101" WHEN "0100100", -- 36
			"00101101000" WHEN "0100101", -- 37
			"00101011001" WHEN "0100110", -- 38
			"00101111000" WHEN "0100111", -- 39

			"00011001101" WHEN "0101000", -- 40
			"00000101011" WHEN "0101001", -- 41
			"00001101011" WHEN "0101010", -- 42
			"01000101011" WHEN "0101011", -- 43

			"00101011010" WHEN "0101100", -- 44
			"01100010000" WHEN "0101101", -- 45
			"00101111001" WHEN "0101110", -- 46
			"01100000000" WHEN "0101111", -- 47

			"00100001101" WHEN "0110000", -- 48
			"00000011100" WHEN "0110001", -- 49
			"00001011100" WHEN "0110010", -- 50
			"01000011100" WHEN "0110011", -- 51

			"00010011100" WHEN "0110100", -- 52
			"01100101000" WHEN "0110101", -- 53
			"00110100001" WHEN "0110110", -- 54
			"01100111000" WHEN "0110111", -- 55

			"00110000011" WHEN "0111000", -- 56
			"00000111011" WHEN "0111001", -- 57
			"00110010001" WHEN "0111010", -- 58
			"00110100000" WHEN "0111011", -- 59

			"00110000010" WHEN "0111100", -- 60
			"00110010000" WHEN "0111101", -- 61
			"00110000001" WHEN "0111110", -- 62
			"00110000000" WHEN "0111111", -- 63

			"00101001101" WHEN "1000000", -- 64
			"00000001110" WHEN "1000001", -- 65
			"00001001110" WHEN "1000010", -- 66
			"00110011000" WHEN "1000011", -- 67

			"00010001110" WHEN "1000100", -- 68
			"00110101000" WHEN "1000101", -- 69
			"00110011001" WHEN "1000110", -- 70
			"00110111000" WHEN "1000111", -- 71

			"00011001110" WHEN "1001000", -- 72
			"10100110000" WHEN "1001001", -- 73
			"00110101001" WHEN "1001010", -- 74
			"10100100000" WHEN "1001011", -- 75

			"00110011010" WHEN "1001100", -- 76
			"10100010000" WHEN "1001101", -- 77
			"00110111001" WHEN "1001110", -- 78
			"10100000000" WHEN "1001111", -- 79

			"00100001110" WHEN "1010000", -- 80
			"00000101100" WHEN "1010001", -- 81
			"00001101100" WHEN "1010010", -- 82
			"01000101100" WHEN "1010011", -- 83

			"00010101100" WHEN "1010100", -- 84
			"10000101100" WHEN "1010101", -- 85
			"01001101100" WHEN "1010110", -- 86
			"10100111000" WHEN "1010111", -- 87

			"00110011011" WHEN "1011000", -- 88
			"01101110000" WHEN "1011001", -- 89
			"01101010001" WHEN "1011010", -- 90
			"01101100000" WHEN "1011011", -- 91

			"00110111010" WHEN "1011100", -- 92
			"01101010000" WHEN "1011101", -- 93
			"01101000001" WHEN "1011110", -- 94
			"01101000000" WHEN "1011111", -- 95

			"00101001110" WHEN "1100000", -- 96
			"00000011101" WHEN "1100001", -- 97
			"00001011101" WHEN "1100010", -- 98
			"01000011101" WHEN "1100011", -- 99

			"00010011101" WHEN "1100100", -- 100
			"01101101000" WHEN "1100101", -- 101
			"01001011101" WHEN "1100110", -- 102
			"01101111000" WHEN "1100111", -- 103

			"00011011101" WHEN "1101000", -- 104
			"11100110000" WHEN "1101001", -- 105
			"01101101001" WHEN "1101010", -- 106
			"11100100000" WHEN "1101011", -- 107

			"00111100010" WHEN "1101100", -- 108
			"11100010000" WHEN "1101101", -- 109
			"01101111001" WHEN "1101110", -- 110
			"11100000000" WHEN "1101111", -- 111

			"00111000100" WHEN "1110000", -- 112
			"00000111100" WHEN "1110001", -- 113
			"00001111100" WHEN "1110010", -- 114
			"01000111100" WHEN "1110011", -- 115

			"00111010010" WHEN "1110100", -- 116
			"10000111100" WHEN "1110101", -- 117
			"00111100001" WHEN "1110110", -- 118
			"11000111100" WHEN "1110111", -- 119

			"00111000011" WHEN "1111000", -- 120
			"00111110000" WHEN "1111001", -- 121
			"00111010001" WHEN "1111010", -- 122
			"00111100000" WHEN "1111011", -- 123

			"00111000010" WHEN "1111100", -- 124
			"00111010000" WHEN "1111101", -- 125
			"00111000001" WHEN "1111110", -- 126
			"00111000000" WHEN "1111111"; -- 127

END behavioral;
